module MaquinaEstados(SW, LEDR, LEDG, KEY);
	input [17:0]SW;
	input [0:0]KEY;
	
	output [17:0]LEDR;
	output [4:0]LEDG;
	
	



endmodule
